module latch_sr(input Set, Reset, Clock
                output Q, Qn);

endmodule